module controle(
	CLOCK, 
	enter,
	reset,
	end_FPGA,
	end_User,
	end_time,
	win,
	match,
	R1,
	R2,
	E1,
	E2,
	E3,
	E4,
	SEL
);

input wire CLOCK, enter, reset, end_FPGA, end_User, end_time, win, match;
output wire R1, R2, E1, E2, E3, E4, SEL;
 
endmodule