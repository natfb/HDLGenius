module Counter_round(

);


endmodule